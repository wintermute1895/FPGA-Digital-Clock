library verilog;
use verilog.vl_types.all;
entity final_test_tb is
end final_test_tb;
