library verilog;
use verilog.vl_types.all;
entity full_functionality_tb is
end full_functionality_tb;
